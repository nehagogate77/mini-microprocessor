LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fsm IS
	PORT (
		clk: IN STD_LOGIC;
		data_in: IN STD_LOGIC;
		reset: IN STD_LOGIC;
		student_id: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		current_state: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE Behavior OF fsm IS
	TYPE state_type IS (s0, s1, s2, s3, s4, s5, s6, s7, s8);
	SIGNAL yfsm: state_type;
	
	BEGIN
		PROCESS(clk, reset)
		BEGIN
			IF reset = '1' THEN
				yfsm <= s0;
			ELSIF (clk'EVENT AND clk = '1') THEN
			CASE yfsm IS
				WHEN s0 =>
					CASE data_in IS
						WHEN '0' => yfsm <= s0;
						WHEN '1' => yfsm <= s1;
					END CASE;
				WHEN s1 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s1;
						WHEN '1' => yfsm <= s2;
					END CASE;
				WHEN s2 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s2;
						WHEN '1' => yfsm <= s3;
					END CASE;
				WHEN s3 =>
					CASE data_in IS
						WHEN '0' => yfsm <= s3;
						WHEN '1' => yfsm <= s4;
					END CASE;
				WHEN s4 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s4;
						WHEN '1' => yfsm <= s5;
					END CASE;
				WHEN s5 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s5;
						WHEN '1' => yfsm <= s6;
					END CASE;
				WHEN s6 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s6;
						WHEN '1' => yfsm <= s7;
					END CASE;
				WHEN s7 =>
					CASE data_in IS
						WHEN '0' => yfsm <= s7;
						WHEN '1' => yfsm <= s8;
					END CASE;
				WHEN s8 => 
					CASE data_in IS
						WHEN '0' => yfsm <= s8;
						WHEN '1' => yfsm <= s0;
					END CASE;
			END CASE;
			END IF;
		END PROCESS;
		PROCESS(yfsm, data_in)
		BEGIN
			CASE yfsm IS
				WHEN s0 => 
					student_id <= "0101";
					current_state <= "0000";
				WHEN s1 => 
					student_id <= "0000";
					current_state <= "0001";
				WHEN s2 => 
					student_id <= "0001";
					current_state <= "0010";
				WHEN s3 => 
					student_id <= "0001";
					current_state <= "0011";
				WHEN s4 => 
					student_id <= "0101";
					current_state <= "0100";
				WHEN s5 => 
					student_id <= "0010";
					current_state <= "0101";
				WHEN s6 => 
					student_id <= "0101";
					current_state <= "0110";
				WHEN s7 => 
					student_id <= "1001";
					current_state <= "0111";
				WHEN s8 => 
					student_id <= "0110";
					current_state <= "1000";
			END CASE;
		END PROCESS;
END Behavior;
